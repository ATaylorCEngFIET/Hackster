
//
// Verific Verilog Description of module lib_pkg
// module not written out since it is a black box. 
//

